//sl2.v
//Coder: Shah-Rukh Khimani
//module designed to shift left logical 2 bits
module shiftLeft2();
	//inputs
	input [3:0] x;
	//outputs
	output [3:0] y;
	//start code
	assign y = x<<2;
//end code
endmodule // end of Module shift left 2
	